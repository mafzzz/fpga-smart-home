module RELAY (input A, input B, output Q);
assign Q = A & B; 
endmodule